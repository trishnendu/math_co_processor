`include "SystemArchHeader.v"

module REG_BANK(
	input wire[`REG_ADDR_WIDTH-1:0] Reg_address
	
	);